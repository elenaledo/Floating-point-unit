module reciprocal(
  input  logic [31:0] data_i,
  output logic [31:0] quoteint,
  output logic []
  output logic [31:0] data_out,
  
);
