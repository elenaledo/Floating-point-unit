module shifter(
  input logic  [7 :0] a_exp_i,
  input logic  [23:0] a_man_i,
  input logic  [7 :0] b_exp_i,
  input logic  [23:0] b_man_i,
  output logic [7 :0] a_exp_o,
  output logic [23:0] a_man_o,
  output logic [7 :0] b_exp_o,
  output logic [23:0] b_man_o,
);

alwa

