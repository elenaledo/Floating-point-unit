module cla(
  input logic [3:0] a,
  input logic [3:0] b,
  input logic       ci,
  output logic[3:0] s,
  output logic      co
);

// p: propagate carry, g: generate carry

  logic [3:0  ] p, g;
always_comb begin
end
